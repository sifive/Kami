Require Export Kami.AllNotations.
(* N.b.: this module exports notations or things dependent on them *)
Require Export Kami.Extraction.
