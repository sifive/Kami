Require Export Kami.AllNoNotations.
(* N.b.: this module exports notations or things dependent on them *)
Require Export Kami.KamiNotations Kami.LibStruct.
Export Word.Notations.
Export ListNotations.
