Require Export AllNoNotations.
(* N.b.: this module exports notations or things dependent on them *)
Require Export KamiNotations LibStruct.
Export Word.Notations.
Export ListNotations.
