Require Export Kami.AllDefn.
(* N.b.: this module exports notations or things dependent on them *)
Require Export Kami.Extraction.
Require Export Kami.Notations Kami.LibStruct.
Export Word.Notations.
Export ListNotations.
